// Header Begin
// Expert list.cdl	19/9/2018
// SINAMICS: Drive
// Header End
r2
p5
p6
p10
p13
p15
r20
r21
r22
r24
r25
r26
r27
r28
r29
r30
r31
r32
r33
r35
r36
r37
r39
p40
p45
r46
r47
r49
r50
r51
r56
r60
r61
r62
r63
r64
r65
r66
r67
r68
r69
r70
r72
r74
r75
r76
r77
r78
r79
r80
r81
r82
r83
r84
r88
r89
r93
r94
p100
r103
p105
r106
r107
r108
r111
p112
p113
r114
p115
r116
p120
p121[0]
p124[0]
p125[0]
r126[0]
r127[0]
r128[0]
p130
p131[0]
p139
p140
p141[0]
p142[0]
p144[0]
p145[0]
r146[0]
r147[0]
r148[0]
p162
p165
r166
p170
p180
p186[0]
r192
p199
r200[0]
p201[0]
r203[0]
r204[0]
r206
r207
r208
r209
p210
p212
r238
p251[0]
p255
p278
p287
r289
p290
r293
p294
p295
r296
r297
p300[0]
p301[0]
r302[0]
r303[0]
p304[0]
p305[0]
p306[0]
p307[0]
p308[0]
p310[0]
p311[0]
r313[0]
p314[0]
p320[0]
p322[0]
p324[0]
p326[0]
r330[0]
r331[0]
r332[0]
r333[0]
p335[0]
r336[0]
r337[0]
r339[0]
p340[0]
p341[0]
p342[0]
p344[0]
p347[0]
p348[0]
p349
p350[0]
p352[0]
p353[0]
p354[0]
p356[0]
p358[0]
p360[0]
p391[0]
p392[0]
p393[0]
r395[0]
r396[0]
p500
p505
p530[0]
p531[0]
p532[0]
p570
p571
p572[0]
p573
p578[0]
p580
p581
p582
p583
r586
r587
r588
r589
p595
p596
p600[0]
p601[0]
p603
p604[0]
p605[0]
p606[0]
p607[0]
p608
p609
p612[0]
p616[0]
p617[0]
p618[0]
p619[0]
p620[0]
p624[0]
p625[0]
p626[0]
p627[0]
p628[0]
p640[0]
p642[0]
p643[0]
p650[0]
p651[0]
p700[0]
p806
r807
p809
p810
p819
p820[0]
p821[0]
p822[0]
p823[0]
p824[0]
p826[0]
p827[0]
p828[0]
r830
p831
r832
p833
r835
r836
r837
r838
p839
p840[0]
p844[0]
p845[0]
p848[0]
p849[0]
p852[0]
p854[0]
p855[0]
p856[0]
p857
p858[0]
p860
p861
p862
r863
p864
p868
p895[0]
r896
p897
r898
r899
p922
r924
p925
r930
r944
r945
r947
r948
r949
p952
p970
p971
r975
r979
p1000[0]
p1001[0]
p1002[0]
p1003[0]
p1004[0]
p1005[0]
p1006[0]
p1007[0]
p1008[0]
p1009[0]
p1010[0]
p1011[0]
p1012[0]
p1013[0]
p1014[0]
p1015[0]
p1020[0]
p1021[0]
p1022[0]
p1023[0]
r1024
p1030[0]
p1035[0]
p1036[0]
p1037[0]
p1038[0]
p1039[0]
p1040[0]
p1041[0]
p1042[0]
p1043[0]
p1044[0]
r1045
p1047[0]
p1048[0]
r1050
p1051[0]
p1052[0]
p1055[0]
p1056[0]
p1058[0]
p1059[0]
p1063[0]
p1070[0]
p1071[0]
r1073
p1075[0]
p1076[0]
r1077
r1078
p1080[0]
p1082[0]
p1083[0]
r1084
p1085[0]
p1086[0]
r1087
p1088[0]
p1091[0]
p1092[0]
p1093[0]
p1094[0]
p1101[0]
p1106[0]
p1110[0]
p1111[0]
r1112
p1113[0]
r1114
p1115
r1119
p1120[0]
p1121[0]
p1122[0]
p1130[0]
p1131[0]
p1134[0]
p1135[0]
p1136[0]
p1137[0]
p1138[0]
p1139[0]
p1140[0]
p1141[0]
p1142[0]
p1143[0]
p1144[0]
p1145[0]
p1148[0]
r1149
r1150
p1151[0]
p1155[0]
p1160[0]
r1169
r1170
p1189[0]
p1190
p1191
p1192[0]
p1193[0]
r1197
r1198
r1199
p1206
p1208
p1210
p1211
p1212
p1213
r1214
p1215
p1216
p1217
p1226[0]
p1227
p1228
p1230[0]
p1231[0]
p1232[0]
p1233[0]
p1234[0]
p1235[0]
p1236[0]
p1237[0]
r1239
p1240[0]
p1244[0]
p1248[0]
p1250[0]
p1278
p1300[0]
p1317[0]
p1318[0]
p1319[0]
p1326[0]
p1327[0]
p1338[0]
p1339[0]
p1345[0]
p1346[0]
p1349[0]
p1400[0]
p1402[0]
p1404[0]
r1406
r1407
r1408
p1409[0]
p1413[0]
p1414[0]
p1415[0]
p1416[0]
p1417[0]
p1418[0]
p1419[0]
p1420[0]
p1421[0]
p1422[0]
p1423[0]
p1424[0]
p1425[0]
p1426[0]
p1428[0]
p1429[0]
p1430[0]
r1432
p1433[0]
p1434[0]
p1435[0]
r1436
r1438
r1439
p1441[0]
r1444
r1445
p1446[0]
p1447[0]
p1448[0]
p1449[0]
p1450[0]
p1451[0]
r1454
p1455[0]
p1456[0]
p1457[0]
p1458[0]
p1459[0]
p1461[0]
p1463[0]
p1464[0]
p1465[0]
p1466[0]
r1468
r1469
p1470[0]
p1472[0]
p1476[0]
p1477[0]
p1478[0]
r1480
r1481
r1482
r1493
p1494[0]
p1497[0]
p1498[0]
p1500[0]
p1501[0]
p1502[0]
r1509
p1511[0]
p1512[0]
p1513[0]
r1515
p1517[0]
r1518
p1520[0]
p1521[0]
p1522[0]
p1523[0]
p1524[0]
p1525[0]
r1526
r1527
p1528[0]
p1529[0]
p1530[0]
p1531[0]
p1532[0]
r1533
r1534
r1535
r1538
r1539
p1542[0]
r1543
p1544
p1545[0]
p1546
r1549
p1550[0]
p1551[0]
p1552[0]
p1554[0]
p1569[0]
p1578[0]
p1579[0]
p1581[0]
p1585[0]
p1590[0]
p1592[0]
p1603[0]
p1612[0]
r1650
r1651
p1656[0]
p1657[0]
p1658[0]
p1659[0]
p1660[0]
p1661[0]
p1662[0]
p1663[0]
p1664[0]
p1665[0]
p1666[0]
p1667[0]
p1668[0]
p1669[0]
p1670[0]
p1671[0]
p1672[0]
p1673[0]
p1674[0]
p1675[0]
p1676[0]
p1699
p1701[0]
p1715[0]
p1717[0]
r1732
r1733
p1755[0]
p1756
r1778
p1780[0]
p1800[0]
p1810
p1815
p1816
p1819
p1821[0]
p1909[0]
p1910
r1912
r1913
r1915
r1927
r1932
r1933
r1934
r1935
r1936
r1937
r1938
r1939
r1947
r1948
r1950
r1951
p1958[0]
p1959[0]
p1960
r1962
r1963
r1969
r1973
p1980[0]
p1981[0]
p1982[0]
p1983
r1984
r1985
r1986
r1987
p1990
p1991[0]
r1992
p1993[0]
p1994[0]
p1995[0]
p1996[0]
p1997[0]
p2000
p2001
p2002
p2003
r2004
p2005
p2006
p2007
r2032
p2037
p2038
p2044
p2045
r2050
p2051
r2053
r2060
p2061
r2063
r2065
r2067
r2074
r2075
r2076
p2079
p2080
p2081
p2082
p2083
p2084
p2088
r2089
r2090
r2091
r2092
r2093
r2094
r2095
p2098
p2099
p2100
p2101
p2103[0]
p2104[0]
p2105[0]
p2106[0]
p2107[0]
p2108[0]
r2109
r2110
p2111
p2112[0]
p2116[0]
p2117[0]
p2118
p2119
r2121
r2122
r2123
r2124
r2125
p2126
p2127
p2128
r2129
r2130
r2131
r2132
r2133
r2134
r2135
r2136
r2138
r2139
p2140[0]
p2141[0]
p2142[0]
p2144[0]
r2145
r2146
p2148[0]
p2149[0]
p2150[0]
p2151[0]
p2153[0]
p2154[0]
p2155[0]
p2156[0]
p2161[0]
p2162[0]
p2163[0]
p2164[0]
p2166[0]
p2167[0]
r2169
p2174[0]
p2175[0]
p2177[0]
p2181[0]
p2182[0]
p2183[0]
p2184[0]
p2185[0]
p2186[0]
p2187[0]
p2188[0]
p2189[0]
p2190[0]
p2192[0]
p2194[0]
p2195[0]
p2196[0]
r2197
r2198
r2199
p2200[0]
p2201[0]
p2202[0]
p2203[0]
p2204[0]
p2205[0]
p2206[0]
p2207[0]
p2208[0]
p2209[0]
p2210[0]
p2211[0]
p2212[0]
p2213[0]
p2214[0]
p2215[0]
p2216[0]
p2220[0]
p2221[0]
p2222[0]
p2223[0]
r2224
r2225
r2229
p2230[0]
r2231
p2235[0]
p2236[0]
p2237[0]
p2238[0]
p2240[0]
r2245
p2247[0]
p2248[0]
r2250
p2252
p2253[0]
p2254[0]
p2255
p2256
p2257
p2258
r2260
p2261
r2262
p2263
p2264[0]
p2265
r2266
p2267
p2268
p2269
p2270
p2271
r2272
r2273
p2274
p2280
p2285
p2286[0]
p2289[0]
p2291
p2292
p2293
r2294
p2295
p2296[0]
p2297[0]
p2298[0]
p2299[0]
p2306
r2349
r2700
r2701
r2702
r2703
r2704
r2705
r2706
r2707
p2810
r2811
p2816
r2817
p2900[0]
p2901[0]
r2902
p2930[0]
p3020
p3041
p3042
p3049[0]
p3050[0]
p3054[0]
p3056[0]
p3058[0]
p3060[0]
p3080
p3081
p3082
p3083
p3088
p3090[0]
p3091[0]
p3092[0]
p3093[0]
p3094[0]
p3095[0]
p3096[0]
p3110
p3111[0]
p3112[0]
r3113
r3115
r3120
r3121
r3122
r3123
r3131
r3132
p3233[0]
p3290
p3291
r3294
p3295
p3296
p3297
p3298
p3299
r3405
p3422
p3510
p3511
p3513
r3517
p3520
p3521
p3523
r3554
p3560
p3562
p3820[0]
p3821[0]
p3822[0]
p3823[0]
p3824[0]
p3825[0]
p3826[0]
p3827[0]
p3828[0]
p3829[0]
p3830[0]
p3831[0]
p3832[0]
p3833[0]
p3834[0]
p3835[0]
p3836[0]
p3837[0]
p3838[0]
p3839[0]
r3840
r3841
p3842
p3845
p3846[0]
p3847[0]
p3870
p3871
p3872
p3873
p3874
r3875
p3876
p3878
p3879
p3900
r3925[0]
r3927[0]
r3928[0]
p3981
p3985
r3986
r3996
r3998[0]
p4600[0]
p4601[0]
p4602[0]
p4603[0]
p4610[0]
p4611[0]
p4612[0]
p4613[0]
r4620
p5007
p5009
r5170
r5171
r5172
r5173
r7760
p7763
p7764[0]
p7770
p8641
p8700
p8701
p8702
p8703
p8704
p8705
p8706
p8707
p8710
p8711
p8712
p8713
p8714
p8715
p8716
p8717
p8720
p8721
p8722
p8723
p8724
p8725
p8726
p8727
p8730
p8731
p8732
p8733
p8734
p8735
p8736
p8737
p8744
r8750
r8751
r8760
r8761
r8784
p8785
p8786
p8787
p8790
r8795
r8796
r8797
p8798
p8837
p8844
r8850
p8851
r8853
r8860
p8861
r8863
r8867
r8874
r8875
r8876
p8880
p8881
p8882
p8883
p8884
p8888
r8889
r8890
r8891
r8892
r8893
r8894
r8895
p8898
p8899
r8960
p9300
p9301
p9302
p9305
p9306
p9307
p9309
p9311
p9312
p9313
p9314
p9315
p9316
p9317
p9318
p9319
p9320
p9321
p9322
p9323
p9324
p9325
p9326
p9328
p9329
p9330
p9331
p9334
p9335
p9341
p9342
p9344
p9345
p9346
p9347
p9348
p9349
p9351
p9352
p9353
p9354
p9355
p9356
p9357
p9358
p9360
p9362
p9363
p9364
p9365
p9366
p9368
p9370
r9371
p9374
p9380
p9381
p9382
p9383
p9385
p9386
p9387
p9388
p9389
r9390
r9398
p9399
r9407
r9408
r9450
r9451
r9490
r9491
r9492
p9493
p9495
p9496
p9497
p9498
p9499
p9500
p9501
p9502
p9505
p9506
p9507
p9509
p9511
p9512
p9513
p9514
p9515
p9516
p9517
p9518
p9519
p9520
p9521
p9522
p9523
p9524
p9525
p9526
p9529
p9530
p9531
p9533
p9534
p9535
p9541
p9542
p9544
p9545
p9546
p9547
p9548
p9549
p9551
p9552
p9553
p9554
p9555
p9556
p9557
p9558
p9559
p9560
p9562
p9563
p9564
p9565
p9566
p9568
p9570
r9571
p9572
p9573
p9574
p9580
p9581
p9582
p9583
p9585
p9586
p9587
p9588
p9589
r9590
p9601
p9602
p9610
p9611
p9620
p9621
p9622
p9650
p9651
p9652
p9653
p9658
p9659
r9660
p9697
p9700
p9701
p9705
r9708
r9710
r9711
r9712
r9713
r9714
r9719
r9720
r9721
r9722
r9723
r9724
r9725
p9726
r9727
r9728
p9729
r9730
r9731
r9732
r9733
r9734
p9740
r9741
r9744
r9745
r9747
r9748
r9749
r9750
p9752
r9753
r9754
r9755
r9756
p9761
p9762
p9763
r9765
r9768
r9769
r9770
r9771
r9772
r9773
r9774
r9780
p9783
r9784
r9785
r9786
r9787
r9794
r9795
r9798
p9799
p9801
p9802
p9810
p9811
p9821
p9822
p9850
p9851
p9852
p9858
r9870
r9871
r9872
r9880
r9881
r9890
r9894
r9895
p9897
r9898
p9899
p60022
